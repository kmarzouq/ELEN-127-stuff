module ROM(addr,data);
	input [9:0]addr;
	reg [11:0]Rt[0:1023];
	output [11:0]data;
	initial begin;
	Rt[0]=0;
	Rt[1]=99;
	Rt[2]=198;
	Rt[3]=297;
	Rt[4]=396;
	Rt[5]=495;
	Rt[6]=594;
	Rt[7]=693;
	Rt[8]=792;
	Rt[9]=891;
	Rt[10]=990;
	Rt[11]=89;
	Rt[12]=188;
	Rt[13]=287;
	Rt[14]=386;
	Rt[15]=485;
	Rt[16]=584;
	Rt[17]=683;
	Rt[18]=782;
	Rt[19]=881;
	Rt[20]=980;
	Rt[21]=79;
	Rt[22]=178;
	Rt[23]=277;
	Rt[24]=376;
	Rt[25]=475;
	Rt[26]=574;
	Rt[27]=673;
	Rt[28]=772;
	Rt[29]=871;
	Rt[30]=970;
	Rt[31]=69;
	Rt[32]=168;
	Rt[33]=267;
	Rt[34]=366;
	Rt[35]=465;
	Rt[36]=564;
	Rt[37]=663;
	Rt[38]=762;
	Rt[39]=861;
	Rt[40]=960;
	Rt[41]=59;
	Rt[42]=158;
	Rt[43]=257;
	Rt[44]=356;
	Rt[45]=455;
	Rt[46]=554;
	Rt[47]=653;
	Rt[48]=752;
	Rt[49]=851;
	Rt[50]=950;
	Rt[51]=49;
	Rt[52]=148;
	Rt[53]=247;
	Rt[54]=346;
	Rt[55]=445;
	Rt[56]=544;
	Rt[57]=643;
	Rt[58]=742;
	Rt[59]=841;
	Rt[60]=940;
	Rt[61]=39;
	Rt[62]=138;
	Rt[63]=237;
	Rt[64]=336;
	Rt[65]=435;
	Rt[66]=534;
	Rt[67]=633;
	Rt[68]=732;
	Rt[69]=831;
	Rt[70]=930;
	Rt[71]=29;
	Rt[72]=128;
	Rt[73]=227;
	Rt[74]=326;
	Rt[75]=425;
	Rt[76]=524;
	Rt[77]=623;
	Rt[78]=722;
	Rt[79]=821;
	Rt[80]=920;
	Rt[81]=19;
	Rt[82]=118;
	Rt[83]=217;
	Rt[84]=316;
	Rt[85]=415;
	Rt[86]=514;
	Rt[87]=613;
	Rt[88]=712;
	Rt[89]=811;
	Rt[90]=910;
	Rt[91]=9;
	Rt[92]=108;
	Rt[93]=207;
	Rt[94]=306;
	Rt[95]=405;
	Rt[96]=504;
	Rt[97]=603;
	Rt[98]=702;
	Rt[99]=801;
	Rt[100]=900;
	Rt[101]=999;
	Rt[102]=98;
	Rt[103]=197;
	Rt[104]=296;
	Rt[105]=395;
	Rt[106]=494;
	Rt[107]=593;
	Rt[108]=692;
	Rt[109]=791;
	Rt[110]=890;
	Rt[111]=989;
	Rt[112]=88;
	Rt[113]=187;
	Rt[114]=286;
	Rt[115]=385;
	Rt[116]=484;
	Rt[117]=583;
	Rt[118]=682;
	Rt[119]=781;
	Rt[120]=880;
	Rt[121]=979;
	Rt[122]=78;
	Rt[123]=177;
	Rt[124]=276;
	Rt[125]=375;
	Rt[126]=474;
	Rt[127]=573;
	Rt[128]=672;
	Rt[129]=771;
	Rt[130]=870;
	Rt[131]=969;
	Rt[132]=68;
	Rt[133]=167;
	Rt[134]=266;
	Rt[135]=365;
	Rt[136]=464;
	Rt[137]=563;
	Rt[138]=662;
	Rt[139]=761;
	Rt[140]=860;
	Rt[141]=959;
	Rt[142]=58;
	Rt[143]=157;
	Rt[144]=256;
	Rt[145]=355;
	Rt[146]=454;
	Rt[147]=553;
	Rt[148]=652;
	Rt[149]=751;
	Rt[150]=850;
	Rt[151]=949;
	Rt[152]=48;
	Rt[153]=147;
	Rt[154]=246;
	Rt[155]=345;
	Rt[156]=444;
	Rt[157]=543;
	Rt[158]=642;
	Rt[159]=741;
	Rt[160]=840;
	Rt[161]=939;
	Rt[162]=38;
	Rt[163]=137;
	Rt[164]=236;
	Rt[165]=335;
	Rt[166]=434;
	Rt[167]=533;
	Rt[168]=632;
	Rt[169]=731;
	Rt[170]=830;
	Rt[171]=929;
	Rt[172]=28;
	Rt[173]=127;
	Rt[174]=226;
	Rt[175]=325;
	Rt[176]=424;
	Rt[177]=523;
	Rt[178]=622;
	Rt[179]=721;
	Rt[180]=820;
	Rt[181]=919;
	Rt[182]=18;
	Rt[183]=117;
	Rt[184]=216;
	Rt[185]=315;
	Rt[186]=414;
	Rt[187]=513;
	Rt[188]=612;
	Rt[189]=711;
	Rt[190]=810;
	Rt[191]=909;
	Rt[192]=8;
	Rt[193]=107;
	Rt[194]=206;
	Rt[195]=305;
	Rt[196]=404;
	Rt[197]=503;
	Rt[198]=602;
	Rt[199]=701;
	Rt[200]=800;
	Rt[201]=899;
	Rt[202]=998;
	Rt[203]=97;
	Rt[204]=196;
	Rt[205]=295;
	Rt[206]=394;
	Rt[207]=493;
	Rt[208]=592;
	Rt[209]=691;
	Rt[210]=790;
	Rt[211]=889;
	Rt[212]=988;
	Rt[213]=87;
	Rt[214]=186;
	Rt[215]=285;
	Rt[216]=384;
	Rt[217]=483;
	Rt[218]=582;
	Rt[219]=681;
	Rt[220]=780;
	Rt[221]=879;
	Rt[222]=978;
	Rt[223]=77;
	Rt[224]=176;
	Rt[225]=275;
	Rt[226]=374;
	Rt[227]=473;
	Rt[228]=572;
	Rt[229]=671;
	Rt[230]=770;
	Rt[231]=869;
	Rt[232]=968;
	Rt[233]=67;
	Rt[234]=166;
	Rt[235]=265;
	Rt[236]=364;
	Rt[237]=463;
	Rt[238]=562;
	Rt[239]=661;
	Rt[240]=760;
	Rt[241]=859;
	Rt[242]=958;
	Rt[243]=57;
	Rt[244]=156;
	Rt[245]=255;
	Rt[246]=354;
	Rt[247]=453;
	Rt[248]=552;
	Rt[249]=651;
	Rt[250]=750;
	Rt[251]=849;
	Rt[252]=948;
	Rt[253]=47;
	Rt[254]=146;
	Rt[255]=245;
	Rt[256]=344;
	Rt[257]=443;
	Rt[258]=542;
	Rt[259]=641;
	Rt[260]=740;
	Rt[261]=839;
	Rt[262]=938;
	Rt[263]=37;
	Rt[264]=136;
	Rt[265]=235;
	Rt[266]=334;
	Rt[267]=433;
	Rt[268]=532;
	Rt[269]=631;
	Rt[270]=730;
	Rt[271]=829;
	Rt[272]=928;
	Rt[273]=27;
	Rt[274]=126;
	Rt[275]=225;
	Rt[276]=324;
	Rt[277]=423;
	Rt[278]=522;
	Rt[279]=621;
	Rt[280]=720;
	Rt[281]=819;
	Rt[282]=918;
	Rt[283]=17;
	Rt[284]=116;
	Rt[285]=215;
	Rt[286]=314;
	Rt[287]=413;
	Rt[288]=512;
	Rt[289]=611;
	Rt[290]=710;
	Rt[291]=809;
	Rt[292]=908;
	Rt[293]=7;
	Rt[294]=106;
	Rt[295]=205;
	Rt[296]=304;
	Rt[297]=403;
	Rt[298]=502;
	Rt[299]=601;
	Rt[300]=700;
	Rt[301]=799;
	Rt[302]=898;
	Rt[303]=997;
	Rt[304]=96;
	Rt[305]=195;
	Rt[306]=294;
	Rt[307]=393;
	Rt[308]=492;
	Rt[309]=591;
	Rt[310]=690;
	Rt[311]=789;
	Rt[312]=888;
	Rt[313]=987;
	Rt[314]=86;
	Rt[315]=185;
	Rt[316]=284;
	Rt[317]=383;
	Rt[318]=482;
	Rt[319]=581;
	Rt[320]=680;
	Rt[321]=779;
	Rt[322]=878;
	Rt[323]=977;
	Rt[324]=76;
	Rt[325]=175;
	Rt[326]=274;
	Rt[327]=373;
	Rt[328]=472;
	Rt[329]=571;
	Rt[330]=670;
	Rt[331]=769;
	Rt[332]=868;
	Rt[333]=967;
	Rt[334]=66;
	Rt[335]=165;
	Rt[336]=264;
	Rt[337]=363;
	Rt[338]=462;
	Rt[339]=561;
	Rt[340]=660;
	Rt[341]=759;
	Rt[342]=858;
	Rt[343]=957;
	Rt[344]=56;
	Rt[345]=155;
	Rt[346]=254;
	Rt[347]=353;
	Rt[348]=452;
	Rt[349]=551;
	Rt[350]=650;
	Rt[351]=749;
	Rt[352]=848;
	Rt[353]=947;
	Rt[354]=46;
	Rt[355]=145;
	Rt[356]=244;
	Rt[357]=343;
	Rt[358]=442;
	Rt[359]=541;
	Rt[360]=640;
	Rt[361]=739;
	Rt[362]=838;
	Rt[363]=937;
	Rt[364]=36;
	Rt[365]=135;
	Rt[366]=234;
	Rt[367]=333;
	Rt[368]=432;
	Rt[369]=531;
	Rt[370]=630;
	Rt[371]=729;
	Rt[372]=828;
	Rt[373]=927;
	Rt[374]=26;
	Rt[375]=125;
	Rt[376]=224;
	Rt[377]=323;
	Rt[378]=422;
	Rt[379]=521;
	Rt[380]=620;
	Rt[381]=719;
	Rt[382]=818;
	Rt[383]=917;
	Rt[384]=16;
	Rt[385]=115;
	Rt[386]=214;
	Rt[387]=313;
	Rt[388]=412;
	Rt[389]=511;
	Rt[390]=610;
	Rt[391]=709;
	Rt[392]=808;
	Rt[393]=907;
	Rt[394]=6;
	Rt[395]=105;
	Rt[396]=204;
	Rt[397]=303;
	Rt[398]=402;
	Rt[399]=501;
	Rt[400]=600;
	Rt[401]=699;
	Rt[402]=798;
	Rt[403]=897;
	Rt[404]=996;
	Rt[405]=95;
	Rt[406]=194;
	Rt[407]=293;
	Rt[408]=392;
	Rt[409]=491;
	Rt[410]=590;
	Rt[411]=689;
	Rt[412]=788;
	Rt[413]=887;
	Rt[414]=986;
	Rt[415]=85;
	Rt[416]=184;
	Rt[417]=283;
	Rt[418]=382;
	Rt[419]=481;
	Rt[420]=580;
	Rt[421]=679;
	Rt[422]=778;
	Rt[423]=877;
	Rt[424]=976;
	Rt[425]=75;
	Rt[426]=174;
	Rt[427]=273;
	Rt[428]=372;
	Rt[429]=471;
	Rt[430]=570;
	Rt[431]=669;
	Rt[432]=768;
	Rt[433]=867;
	Rt[434]=966;
	Rt[435]=65;
	Rt[436]=164;
	Rt[437]=263;
	Rt[438]=362;
	Rt[439]=461;
	Rt[440]=560;
	Rt[441]=659;
	Rt[442]=758;
	Rt[443]=857;
	Rt[444]=956;
	Rt[445]=55;
	Rt[446]=154;
	Rt[447]=253;
	Rt[448]=352;
	Rt[449]=451;
	Rt[450]=550;
	Rt[451]=649;
	Rt[452]=748;
	Rt[453]=847;
	Rt[454]=946;
	Rt[455]=45;
	Rt[456]=144;
	Rt[457]=243;
	Rt[458]=342;
	Rt[459]=441;
	Rt[460]=540;
	Rt[461]=639;
	Rt[462]=738;
	Rt[463]=837;
	Rt[464]=936;
	Rt[465]=35;
	Rt[466]=134;
	Rt[467]=233;
	Rt[468]=332;
	Rt[469]=431;
	Rt[470]=530;
	Rt[471]=629;
	Rt[472]=728;
	Rt[473]=827;
	Rt[474]=926;
	Rt[475]=25;
	Rt[476]=124;
	Rt[477]=223;
	Rt[478]=322;
	Rt[479]=421;
	Rt[480]=520;
	Rt[481]=619;
	Rt[482]=718;
	Rt[483]=817;
	Rt[484]=916;
	Rt[485]=15;
	Rt[486]=114;
	Rt[487]=213;
	Rt[488]=312;
	Rt[489]=411;
	Rt[490]=510;
	Rt[491]=609;
	Rt[492]=708;
	Rt[493]=807;
	Rt[494]=906;
	Rt[495]=5;
	Rt[496]=104;
	Rt[497]=203;
	Rt[498]=302;
	Rt[499]=401;
	Rt[500]=500;
	Rt[501]=599;
	Rt[502]=698;
	Rt[503]=797;
	Rt[504]=896;
	Rt[505]=995;
	Rt[506]=94;
	Rt[507]=193;
	Rt[508]=292;
	Rt[509]=391;
	Rt[510]=490;
	Rt[511]=589;
	Rt[512]=688;
	Rt[513]=787;
	Rt[514]=886;
	Rt[515]=985;
	Rt[516]=84;
	Rt[517]=183;
	Rt[518]=282;
	Rt[519]=381;
	Rt[520]=480;
	Rt[521]=579;
	Rt[522]=678;
	Rt[523]=777;
	Rt[524]=876;
	Rt[525]=975;
	Rt[526]=74;
	Rt[527]=173;
	Rt[528]=272;
	Rt[529]=371;
	Rt[530]=470;
	Rt[531]=569;
	Rt[532]=668;
	Rt[533]=767;
	Rt[534]=866;
	Rt[535]=965;
	Rt[536]=64;
	Rt[537]=163;
	Rt[538]=262;
	Rt[539]=361;
	Rt[540]=460;
	Rt[541]=559;
	Rt[542]=658;
	Rt[543]=757;
	Rt[544]=856;
	Rt[545]=955;
	Rt[546]=54;
	Rt[547]=153;
	Rt[548]=252;
	Rt[549]=351;
	Rt[550]=450;
	Rt[551]=549;
	Rt[552]=648;
	Rt[553]=747;
	Rt[554]=846;
	Rt[555]=945;
	Rt[556]=44;
	Rt[557]=143;
	Rt[558]=242;
	Rt[559]=341;
	Rt[560]=440;
	Rt[561]=539;
	Rt[562]=638;
	Rt[563]=737;
	Rt[564]=836;
	Rt[565]=935;
	Rt[566]=34;
	Rt[567]=133;
	Rt[568]=232;
	Rt[569]=331;
	Rt[570]=430;
	Rt[571]=529;
	Rt[572]=628;
	Rt[573]=727;
	Rt[574]=826;
	Rt[575]=925;
	Rt[576]=24;
	Rt[577]=123;
	Rt[578]=222;
	Rt[579]=321;
	Rt[580]=420;
	Rt[581]=519;
	Rt[582]=618;
	Rt[583]=717;
	Rt[584]=816;
	Rt[585]=915;
	Rt[586]=14;
	Rt[587]=113;
	Rt[588]=212;
	Rt[589]=311;
	Rt[590]=410;
	Rt[591]=509;
	Rt[592]=608;
	Rt[593]=707;
	Rt[594]=806;
	Rt[595]=905;
	Rt[596]=4;
	Rt[597]=103;
	Rt[598]=202;
	Rt[599]=301;
	Rt[600]=400;
	Rt[601]=499;
	Rt[602]=598;
	Rt[603]=697;
	Rt[604]=796;
	Rt[605]=895;
	Rt[606]=994;
	Rt[607]=93;
	Rt[608]=192;
	Rt[609]=291;
	Rt[610]=390;
	Rt[611]=489;
	Rt[612]=588;
	Rt[613]=687;
	Rt[614]=786;
	Rt[615]=885;
	Rt[616]=984;
	Rt[617]=83;
	Rt[618]=182;
	Rt[619]=281;
	Rt[620]=380;
	Rt[621]=479;
	Rt[622]=578;
	Rt[623]=677;
	Rt[624]=776;
	Rt[625]=875;
	Rt[626]=974;
	Rt[627]=73;
	Rt[628]=172;
	Rt[629]=271;
	Rt[630]=370;
	Rt[631]=469;
	Rt[632]=568;
	Rt[633]=667;
	Rt[634]=766;
	Rt[635]=865;
	Rt[636]=964;
	Rt[637]=63;
	Rt[638]=162;
	Rt[639]=261;
	Rt[640]=360;
	Rt[641]=459;
	Rt[642]=558;
	Rt[643]=657;
	Rt[644]=756;
	Rt[645]=855;
	Rt[646]=954;
	Rt[647]=53;
	Rt[648]=152;
	Rt[649]=251;
	Rt[650]=350;
	Rt[651]=449;
	Rt[652]=548;
	Rt[653]=647;
	Rt[654]=746;
	Rt[655]=845;
	Rt[656]=944;
	Rt[657]=43;
	Rt[658]=142;
	Rt[659]=241;
	Rt[660]=340;
	Rt[661]=439;
	Rt[662]=538;
	Rt[663]=637;
	Rt[664]=736;
	Rt[665]=835;
	Rt[666]=934;
	Rt[667]=33;
	Rt[668]=132;
	Rt[669]=231;
	Rt[670]=330;
	Rt[671]=429;
	Rt[672]=528;
	Rt[673]=627;
	Rt[674]=726;
	Rt[675]=825;
	Rt[676]=924;
	Rt[677]=23;
	Rt[678]=122;
	Rt[679]=221;
	Rt[680]=320;
	Rt[681]=419;
	Rt[682]=518;
	Rt[683]=617;
	Rt[684]=716;
	Rt[685]=815;
	Rt[686]=914;
	Rt[687]=13;
	Rt[688]=112;
	Rt[689]=211;
	Rt[690]=310;
	Rt[691]=409;
	Rt[692]=508;
	Rt[693]=607;
	Rt[694]=706;
	Rt[695]=805;
	Rt[696]=904;
	Rt[697]=3;
	Rt[698]=102;
	Rt[699]=201;
	Rt[700]=300;
	Rt[701]=399;
	Rt[702]=498;
	Rt[703]=597;
	Rt[704]=696;
	Rt[705]=795;
	Rt[706]=894;
	Rt[707]=993;
	Rt[708]=92;
	Rt[709]=191;
	Rt[710]=290;
	Rt[711]=389;
	Rt[712]=488;
	Rt[713]=587;
	Rt[714]=686;
	Rt[715]=785;
	Rt[716]=884;
	Rt[717]=983;
	Rt[718]=82;
	Rt[719]=181;
	Rt[720]=280;
	Rt[721]=379;
	Rt[722]=478;
	Rt[723]=577;
	Rt[724]=676;
	Rt[725]=775;
	Rt[726]=874;
	Rt[727]=973;
	Rt[728]=72;
	Rt[729]=171;
	Rt[730]=270;
	Rt[731]=369;
	Rt[732]=468;
	Rt[733]=567;
	Rt[734]=666;
	Rt[735]=765;
	Rt[736]=864;
	Rt[737]=963;
	Rt[738]=62;
	Rt[739]=161;
	Rt[740]=260;
	Rt[741]=359;
	Rt[742]=458;
	Rt[743]=557;
	Rt[744]=656;
	Rt[745]=755;
	Rt[746]=854;
	Rt[747]=953;
	Rt[748]=52;
	Rt[749]=151;
	Rt[750]=250;
	Rt[751]=349;
	Rt[752]=448;
	Rt[753]=547;
	Rt[754]=646;
	Rt[755]=745;
	Rt[756]=844;
	Rt[757]=943;
	Rt[758]=42;
	Rt[759]=141;
	Rt[760]=240;
	Rt[761]=339;
	Rt[762]=438;
	Rt[763]=537;
	Rt[764]=636;
	Rt[765]=735;
	Rt[766]=834;
	Rt[767]=933;
	Rt[768]=32;
	Rt[769]=131;
	Rt[770]=230;
	Rt[771]=329;
	Rt[772]=428;
	Rt[773]=527;
	Rt[774]=626;
	Rt[775]=725;
	Rt[776]=824;
	Rt[777]=923;
	Rt[778]=22;
	Rt[779]=121;
	Rt[780]=220;
	Rt[781]=319;
	Rt[782]=418;
	Rt[783]=517;
	Rt[784]=616;
	Rt[785]=715;
	Rt[786]=814;
	Rt[787]=913;
	Rt[788]=12;
	Rt[789]=111;
	Rt[790]=210;
	Rt[791]=309;
	Rt[792]=408;
	Rt[793]=507;
	Rt[794]=606;
	Rt[795]=705;
	Rt[796]=804;
	Rt[797]=903;
	Rt[798]=2;
	Rt[799]=101;
	Rt[800]=200;
	Rt[801]=299;
	Rt[802]=398;
	Rt[803]=497;
	Rt[804]=596;
	Rt[805]=695;
	Rt[806]=794;
	Rt[807]=893;
	Rt[808]=992;
	Rt[809]=91;
	Rt[810]=190;
	Rt[811]=289;
	Rt[812]=388;
	Rt[813]=487;
	Rt[814]=586;
	Rt[815]=685;
	Rt[816]=784;
	Rt[817]=883;
	Rt[818]=982;
	Rt[819]=81;
	Rt[820]=180;
	Rt[821]=279;
	Rt[822]=378;
	Rt[823]=477;
	Rt[824]=576;
	Rt[825]=675;
	Rt[826]=774;
	Rt[827]=873;
	Rt[828]=972;
	Rt[829]=71;
	Rt[830]=170;
	Rt[831]=269;
	Rt[832]=368;
	Rt[833]=467;
	Rt[834]=566;
	Rt[835]=665;
	Rt[836]=764;
	Rt[837]=863;
	Rt[838]=962;
	Rt[839]=61;
	Rt[840]=160;
	Rt[841]=259;
	Rt[842]=358;
	Rt[843]=457;
	Rt[844]=556;
	Rt[845]=655;
	Rt[846]=754;
	Rt[847]=853;
	Rt[848]=952;
	Rt[849]=51;
	Rt[850]=150;
	Rt[851]=249;
	Rt[852]=348;
	Rt[853]=447;
	Rt[854]=546;
	Rt[855]=645;
	Rt[856]=744;
	Rt[857]=843;
	Rt[858]=942;
	Rt[859]=41;
	Rt[860]=140;
	Rt[861]=239;
	Rt[862]=338;
	Rt[863]=437;
	Rt[864]=536;
	Rt[865]=635;
	Rt[866]=734;
	Rt[867]=833;
	Rt[868]=932;
	Rt[869]=31;
	Rt[870]=130;
	Rt[871]=229;
	Rt[872]=328;
	Rt[873]=427;
	Rt[874]=526;
	Rt[875]=625;
	Rt[876]=724;
	Rt[877]=823;
	Rt[878]=922;
	Rt[879]=21;
	Rt[880]=120;
	Rt[881]=219;
	Rt[882]=318;
	Rt[883]=417;
	Rt[884]=516;
	Rt[885]=615;
	Rt[886]=714;
	Rt[887]=813;
	Rt[888]=912;
	Rt[889]=11;
	Rt[890]=110;
	Rt[891]=209;
	Rt[892]=308;
	Rt[893]=407;
	Rt[894]=506;
	Rt[895]=605;
	Rt[896]=704;
	Rt[897]=803;
	Rt[898]=902;
	Rt[899]=1;
	Rt[900]=100;
	Rt[901]=199;
	Rt[902]=298;
	Rt[903]=397;
	Rt[904]=496;
	Rt[905]=595;
	Rt[906]=694;
	Rt[907]=793;
	Rt[908]=892;
	Rt[909]=991;
	Rt[910]=90;
	Rt[911]=189;
	Rt[912]=288;
	Rt[913]=387;
	Rt[914]=486;
	Rt[915]=585;
	Rt[916]=684;
	Rt[917]=783;
	Rt[918]=882;
	Rt[919]=981;
	Rt[920]=80;
	Rt[921]=179;
	Rt[922]=278;
	Rt[923]=377;
	Rt[924]=476;
	Rt[925]=575;
	Rt[926]=674;
	Rt[927]=773;
	Rt[928]=872;
	Rt[929]=971;
	Rt[930]=70;
	Rt[931]=169;
	Rt[932]=268;
	Rt[933]=367;
	Rt[934]=466;
	Rt[935]=565;
	Rt[936]=664;
	Rt[937]=763;
	Rt[938]=862;
	Rt[939]=961;
	Rt[940]=60;
	Rt[941]=159;
	Rt[942]=258;
	Rt[943]=357;
	Rt[944]=456;
	Rt[945]=555;
	Rt[946]=654;
	Rt[947]=753;
	Rt[948]=852;
	Rt[949]=951;
	Rt[950]=50;
	Rt[951]=149;
	Rt[952]=248;
	Rt[953]=347;
	Rt[954]=446;
	Rt[955]=545;
	Rt[956]=644;
	Rt[957]=743;
	Rt[958]=842;
	Rt[959]=941;
	Rt[960]=40;
	Rt[961]=139;
	Rt[962]=238;
	Rt[963]=337;
	Rt[964]=436;
	Rt[965]=535;
	Rt[966]=634;
	Rt[967]=733;
	Rt[968]=832;
	Rt[969]=931;
	Rt[970]=30;
	Rt[971]=129;
	Rt[972]=228;
	Rt[973]=327;
	Rt[974]=426;
	Rt[975]=525;
	Rt[976]=624;
	Rt[977]=723;
	Rt[978]=822;
	Rt[979]=921;
	Rt[980]=20;
	Rt[981]=119;
	Rt[982]=218;
	Rt[983]=317;
	Rt[984]=416;
	Rt[985]=515;
	Rt[986]=614;
	Rt[987]=713;
	Rt[988]=812;
	Rt[989]=911;
	Rt[990]=10;
	Rt[991]=109;
	Rt[992]=208;
	Rt[993]=307;
	Rt[994]=406;
	Rt[995]=505;
	Rt[996]=604;
	Rt[997]=703;
	Rt[998]=802;
	Rt[999]=901;
	Rt[1000]=0;
	Rt[1001]=99;
	Rt[1002]=198;
	Rt[1003]=297;
	Rt[1004]=396;
	Rt[1005]=495;
	Rt[1006]=594;
	Rt[1007]=693;
	Rt[1008]=792;
	Rt[1009]=891;
	Rt[1010]=990;
	Rt[1011]=89;
	Rt[1012]=188;
	Rt[1013]=287;
	Rt[1014]=386;
	Rt[1015]=485;
	Rt[1016]=584;
	Rt[1017]=683;
	Rt[1018]=782;
	Rt[1019]=881;
	Rt[1020]=980;
	Rt[1021]=79;
	Rt[1022]=178;
	Rt[1023]=277;
	end;
	assign data = Rt[addr]; 
 endmodule